`timescale 1ns / 1ps

module SpartanBreakout(
   input CLK_50M,
   output AUDIO_OUT
   );

   AudioPlayer player(.CLK(CLK_50M), .AUDIO(AUDIO_OUT));
endmodule
